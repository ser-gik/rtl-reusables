
`ifndef REUSABLES_VH
`define REUSABLES_VH

`define R_STATIC_ERROR(msg) msg err()

`endif

