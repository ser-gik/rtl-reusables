
`ifndef UART_8N1
`define UART_8N1

`define UART_8N1_BAUD_9600 2'b01
`define UART_8N1_BAUD_19200 2'b10

`endif // UART_8N1
